
localparam ALU_AND = 4'b0000;
localparam ALU_OR  = 4'b0001;
localparam ALU_ADD = 4'b0010;
localparam ALU_SUB = 4'b0110;
localparam ALU_EQ  = 4'b0111;
localparam ALU_NOP = 4'b1111;
