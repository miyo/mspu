
/******************************************************
 * ALU OP
 ******************************************************/
localparam ALU_AND = 4'b0000;
localparam ALU_OR  = 4'b0001;
localparam ALU_XOR = 4'b0010;
localparam ALU_ADD = 4'b0100;
localparam ALU_SUB = 4'b0101;
localparam ALU_EQ  = 4'b1000;
localparam ALU_NE  = 4'b1001;
localparam ALU_LT  = 4'b1010;
localparam ALU_GE  = 4'b1011;

/******************************************************
 * MUL OP
 ******************************************************/
localparam MUL_NOP    = 4'b0000;
localparam MUL_MUL    = 4'b0001;
localparam MUL_MULH   = 4'b0010;
localparam MUL_MULHSU = 4'b0011;
localparam MUL_MULHU  = 4'b0100;

/******************************************************
 * ISA
 ******************************************************/

// RV32I
localparam LUI   = 32'b????????????????????_?????_0110111;
localparam AUIPC = 32'b????????????????????_?????_0010111;

localparam JAL   = 32'b????????????????????_?????_1101111;
localparam JALR  = 32'b????????????_?????_000_?????_1100111;

localparam BEQ   = 32'b???????_?????_?????_000_?????_1100011;
localparam BNE   = 32'b???????_?????_?????_001_?????_1100011;
localparam BLT   = 32'b???????_?????_?????_100_?????_1100011;
localparam BGE   = 32'b???????_?????_?????_101_?????_1100011;
localparam BLTU  = 32'b???????_?????_?????_110_?????_1100011;
localparam BGEU  = 32'b???????_?????_?????_111_?????_1100011;

localparam LB    = 32'b????????????_?????_000_?????_0000011;
localparam LH    = 32'b????????????_?????_001_?????_0000011;
localparam LW    = 32'b????????????_?????_010_?????_0000011;
localparam LBU   = 32'b????????????_?????_100_?????_0000011;
localparam LHU   = 32'b????????????_?????_101_?????_0000011;

localparam SB    = 32'b???????_?????_?????_000_?????_0100011;
localparam SH    = 32'b???????_?????_?????_001_?????_0100011;
localparam SW    = 32'b???????_?????_?????_010_?????_0100011;

localparam ADDI  = 32'b????????????_?????_000_?????_0010011;
localparam SLTI  = 32'b????????????_?????_010_?????_0010011;
localparam SLTIU = 32'b????????????_?????_011_?????_0010011;
localparam XORI  = 32'b????????????_?????_100_?????_0010011;
localparam ORI   = 32'b????????????_?????_110_?????_0010011;
localparam ANDI  = 32'b????????????_?????_111_?????_0010011;

localparam SLLI  = 32'b0000000_?????_?????_001_?????_0010011;
localparam SRLI  = 32'b0000000_?????_?????_101_?????_0010011;
localparam SRAI  = 32'b0100000_?????_?????_101_?????_0010011;

localparam ADD   = 32'b0000000_?????_?????_000_?????_0110011;
localparam SUB   = 32'b0100000_?????_?????_000_?????_0110011;
localparam SLL   = 32'b0000000_?????_?????_001_?????_0110011;
localparam SLT   = 32'b0000000_?????_?????_010_?????_0110011;
localparam SLTU  = 32'b0000000_?????_?????_011_?????_0110011;
localparam XOR   = 32'b0000000_?????_?????_100_?????_0110011;
localparam SRL   = 32'b0000000_?????_?????_101_?????_0110011;
localparam SRA   = 32'b0100000_?????_?????_101_?????_0110011;
localparam OR    = 32'b0000000_?????_?????_110_?????_0110011;
localparam AND   = 32'b0100000_?????_?????_111_?????_0110011;

localparam FENCE   = 32'b0000_????_????_00000_000_00000_0001111;
localparam FENCE_I = 32'b0000_0000_0000_00000_001_00000_0001111;

localparam ECALL  = 32'b000000000000_00000_000_00000_1110011;
localparam EBREAK = 32'b000000000001_00000_000_00000_1110011;

localparam CSRRW  = 32'b????????????_?????_001_?????_1110011;
localparam CSRRS  = 32'b????????????_?????_010_?????_1110011;
localparam CSRRC  = 32'b????????????_?????_011_?????_1110011;
localparam CSRRWI = 32'b????????????_?????_101_?????_1110011;
localparam CSRRSI = 32'b????????????_?????_110_?????_1110011;
localparam CSRRCI = 32'b????????????_?????_111_?????_1110011;

// RV64I
localparam LWU = 32'b????????????_?????_110_?????_0000011;
localparam LD  = 32'b????????????_?????_011_?????_0000011;

localparam SD  = 32'b???????_?????_?????_011_?????_0100011;

localparam ADDIW = 32'b????????????_?????_000_?????_0011011;
localparam SLLIW = 32'b0000000_?????_?????_001_?????_0011011;
localparam SRLIW = 32'b0000000_?????_?????_101_?????_0011011;
localparam SRAIW = 32'b0100000_?????_?????_101_?????_0011011;

localparam ADDW = 32'b0000000_?????_?????_000_?????_0111011;
localparam SUBW = 32'b0100000_?????_?????_000_?????_0111011;
localparam SLLW = 32'b0000000_?????_?????_001_?????_0111011;
localparam SRLW = 32'b0000000_?????_?????_101_?????_0111011;
localparam SRAW = 32'b0100000_?????_?????_101_?????_0111011;

// RV32M
localparam MUL    = 32'b0000001_?????_?????_000_?????_0110011;
localparam MULH   = 32'b0000001_?????_?????_001_?????_0110011;
localparam MULHSU = 32'b0000001_?????_?????_010_?????_0110011;
localparam MULHU  = 32'b0000001_?????_?????_011_?????_0110011;
localparam DIV    = 32'b0000001_?????_?????_100_?????_0110011;
localparam DIVU   = 32'b0000001_?????_?????_101_?????_0110011;
localparam REM    = 32'b0000001_?????_?????_110_?????_0110011;
localparam REMU   = 32'b0000001_?????_?????_111_?????_0110011;

// RV64M
localparam MULW  = 32'b0000001_?????_?????_000_?????_0111011;
localparam DIVW  = 32'b0000001_?????_?????_100_?????_0111011;
localparam DIVUW = 32'b0000001_?????_?????_101_?????_0111011;
localparam REMW  = 32'b0000001_?????_?????_110_?????_0111011;
localparam REMUW = 32'b0000001_?????_?????_111_?????_0111011;

// RV32A
localparam LR_W      = 32'b00010_?_?_00000_?????_010_?????_0101111;
localparam SC_W      = 32'b00011_?_?_?????_?????_010_?????_0101111;
localparam AMOSWAP_W = 32'b00001_?_?_?????_?????_010_?????_0101111;
localparam AMOADD_W  = 32'b00000_?_?_?????_?????_010_?????_0101111;
localparam AMOXOR_W  = 32'b00100_?_?_?????_?????_010_?????_0101111;
localparam AMOAND_W  = 32'b01100_?_?_?????_?????_010_?????_0101111;
localparam AMOOR_W   = 32'b01000_?_?_?????_?????_010_?????_0101111;
localparam AMOMIN_W  = 32'b10000_?_?_?????_?????_010_?????_0101111;
localparam AMOMAX_W  = 32'b10100_?_?_?????_?????_010_?????_0101111;
localparam AMOMINU_W = 32'b11000_?_?_?????_?????_010_?????_0101111;
localparam AMOMAXU_W = 32'b11100_?_?_?????_?????_010_?????_0101111;

// RV64A
localparam LR_D      = 32'b00010_?_?_00000_?????_011_?????_0101111;
localparam SC_D      = 32'b00011_?_?_?????_?????_011_?????_0101111;
localparam AMOSWAP_D = 32'b00001_?_?_?????_?????_011_?????_0101111;
localparam AMOADD_D  = 32'b00000_?_?_?????_?????_011_?????_0101111;
localparam AMOXOR_D  = 32'b00100_?_?_?????_?????_011_?????_0101111;
localparam AMOAND_D  = 32'b01100_?_?_?????_?????_011_?????_0101111;
localparam AMOOR_D   = 32'b01000_?_?_?????_?????_011_?????_0101111;
localparam AMOMIN_D  = 32'b10000_?_?_?????_?????_011_?????_0101111;
localparam AMOMAX_D  = 32'b10100_?_?_?????_?????_011_?????_0101111;
localparam AMOMINU_D = 32'b11000_?_?_?????_?????_011_?????_0101111;
localparam AMOMAXU_D = 32'b11100_?_?_?????_?????_011_?????_0101111;

// RV32F
localparam FLW = 32'b????????????_?????_010_?????_0000111;
localparam FSW = 32'b???????_?????_?????_010_?????_0100111;

localparam FMADD_S  = 32'b?????_00_?????_?????_???_?????_1000011;
localparam FMSUB_S  = 32'b?????_00_?????_?????_???_?????_1000111;
localparam FNMSUB_S = 32'b?????_00_?????_?????_???_?????_1001011;
localparam FNMADD_S = 32'b?????_00_?????_?????_???_?????_1001111;

localparam FADD_S    = 32'b0000000_?????_?????_???_?????_1010011;
localparam FSUB_S    = 32'b0000100_?????_?????_???_?????_1010011;
localparam FMUL_S    = 32'b0001000_?????_?????_???_?????_1010011;
localparam FDIV_S    = 32'b0001100_?????_?????_???_?????_1010011;
localparam FSQRT_S   = 32'b0101100_00000_?????_???_?????_1010011;
localparam FSGNJ_S   = 32'b0010000_?????_?????_000_?????_1010011;
localparam FSGNJN_S  = 32'b0010000_?????_?????_001_?????_1010011;
localparam FSGNJX_S  = 32'b0010000_?????_?????_010_?????_1010011;
localparam FMIN_S    = 32'b0010100_?????_?????_000_?????_1010011;
localparam FMAX_S    = 32'b0010100_?????_?????_001_?????_1010011;
localparam FCVT_W_S  = 32'b1100000_00000_?????_???_?????_1010011;
localparam FCVT_WU_S = 32'b1100000_00001_?????_???_?????_1010011;
localparam FMV_X_W   = 32'b1110000_00000_?????_000_?????_1010011;
localparam FEQ_S     = 32'b1010000_?????_?????_010_?????_1010011;
localparam FLT_S     = 32'b1010000_?????_?????_001_?????_1010011;
localparam FLE_S     = 32'b1010000_?????_?????_000_?????_1010011;
localparam FCLASS_S  = 32'b1110000_00000_?????_001_?????_1010011;
localparam FCVT_S_W  = 32'b1101000_00000_?????_???_?????_1010011;
localparam FCVT_S_WU = 32'b1101000_00001_?????_???_?????_1010011;
localparam FMV_W_X   = 32'b1111000_00000_?????_000_?????_1010011;

// RV64F
localparam FCVT_L_S  = 32'b1100000_00010_?????_???_?????_1010011;
localparam FCVT_LU_S = 32'b1100000_00011_?????_???_?????_1010011;
localparam FCVT_S_L  = 32'b1101000_00010_?????_???_?????_1010011;
localparam FCVT_S_LU = 32'b1101000_00011_?????_???_?????_1010011;

// RV32D
localparam FLD = 32'b????????????_?????_011_?????_0000111;
localparam FSD = 32'b???????_?????_?????_011_?????_0100111;

localparam FMADD_D  = 32'b?????_01_?????_?????_???_?????_1000011;
localparam FMSUB_D  = 32'b?????_01_?????_?????_???_?????_1000111;
localparam FNMSUB_D = 32'b?????_01_?????_?????_???_?????_1001011;
localparam FNMADD_D = 32'b?????_01_?????_?????_???_?????_1001111;

localparam FADD_D    = 32'b0000001_?????_?????_???_?????_1010011;
localparam FSUB_D    = 32'b0000101_?????_?????_???_?????_1010011;
localparam FMUL_D    = 32'b0001001_?????_?????_???_?????_1010011;
localparam FDIV_D    = 32'b0001101_?????_?????_???_?????_1010011;
localparam FSQRT_D   = 32'b0101101_00000_?????_???_?????_1010011;
localparam FSGNJ_D   = 32'b0010001_?????_?????_000_?????_1010011;
localparam FSGNJN_D  = 32'b0010001_?????_?????_001_?????_1010011;
localparam FSGNJX_D  = 32'b0010001_?????_?????_010_?????_1010011;
localparam FMIN_D    = 32'b0010101_?????_?????_000_?????_1010011;
localparam FMAX_D    = 32'b0010101_?????_?????_001_?????_1010011;
localparam FCVT_S_D  = 32'b0100000_00001_?????_???_?????_1010011;
localparam FCVT_D_S  = 32'b0100001_00000_?????_???_?????_1010011;
localparam FEQ_D     = 32'b1010001_?????_?????_010_?????_1010011;
localparam FLT_D     = 32'b1010001_?????_?????_001_?????_1010011;
localparam FLE_D     = 32'b1010001_?????_?????_000_?????_1010011;
localparam FCLASS_D  = 32'b1110001_00000_?????_001_?????_1010011;
localparam FCVT_W_D  = 32'b1100001_00000_?????_???_?????_1010011;
localparam FCVT_WU_D = 32'b1100001_00001_?????_???_?????_1010011;
localparam FCVT_D_W  = 32'b1101001_00000_?????_???_?????_1010011;
localparam FCVT_D_WU = 32'b1101001_00001_?????_???_?????_1010011;

// RV64D
localparam FCVT_L_D  = 32'b1100001_00010_?????_???_?????_1010011;
localparam FCVT_LU_D = 32'b1100001_00011_?????_???_?????_1010011;
localparam FMV_X_D   = 32'b1110001_00000_?????_000_?????_1010011;
localparam FCVT_D_L  = 32'b1101001_00010_?????_???_?????_1010011;
localparam FCVT_D_LU = 32'b1101001_00011_?????_???_?????_1010011;
localparam FMV_D_X   = 32'b1111001_00000_?????_000_?????_1010011;
